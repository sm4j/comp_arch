--Data Flip Flop Positive-Edge Triggered
--Behavioral Model
--Jordan Small, Nov. 4, 2023

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY DFF_SmallJordan IS
PORT (
		D, Clock : IN    STD_LOGIC;
		   Q, QN : INOUT STD_LOGIC
	 );
END DFF_SmallJordan;

ARCHITECTURE behavior OF DFF_SmallJordan IS
BEGIN
--Update register output on the clock's rising edge
	PROCESS (Clock)
	BEGIN
		IF (rising_edge(clock)) THEN
			Q <= D;
		END IF;
	END PROCESS;
END behavior;